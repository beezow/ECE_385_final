module centroid
(	
input logic image[307200],
output logic[10:0] x,y
);

always_comb begin





end

endmodule