//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Viral Mehta                                                        --
//    Spring 2005                                                        --
//                                                                       --
//    Modified by Stephen Kempf 03-01-2006                               --
//                              03-12-2007                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 298 Lab 7                                         --
//    UIUC ECE Department                                                --
//-------------------------------------------------------------------------
module  ball ( input Reset, frame_clk,
					input [9:0] PaddleX, PaddleY, PaddleS,
					output [3:0] Score1, Score2,
               output [9:0]  BallX, BallY, BallS);
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion, Ball_Size;
	 
    parameter [9:0] Ball_X_Center=320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center=240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min=0;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max=639;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min=0;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max=479;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step=3;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step=3;      // Step size on the Y axis

    assign Ball_Size = 4;  // assigns the value 4 as a 10-digit binary number, ie "0000000100"

    int DistX, DistY;
	 assign DistX = PaddleX - Ball_X_Pos;
    assign DistY = PaddleY - Ball_Y_Pos;

	 logic in_paddle;
	 assign in_paddle = ((DistX*DistX/8) + ( DistY*DistY/(PaddleS*PaddleS) ) <= 1);
		
    always_ff @ (posedge Reset or posedge frame_clk )
    begin: Move_Ball
        if (Reset)  // Asynchronous Reset
        begin 
           // Ball_Y_Motion <= 10'd0; //Ball_Y_Step;
			//	Ball_X_Motion <= 10'd0; //Ball_X_Step;
				Ball_Y_Pos <= Ball_Y_Center;
				Ball_X_Pos <= Ball_X_Center;
				
				Ball_X_Motion <= 3;//A
				Ball_Y_Motion <= -3;
				Score1 <=0;
				Score2 <=0;

        end
           
        else 
        begin 
				 if (Score1<=9 && Score2<=9) begin 
					 if ( (Ball_Y_Pos + Ball_Size-1) >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
						  Ball_Y_Motion <= (~ (Ball_Y_Step) + 1'b1);  // 2's complement.
						  
					 else if ( (Ball_Y_Pos - Ball_Size+1) <= Ball_Y_Min )  // Ball is at the top edge, BOUNCE!
						  Ball_Y_Motion <= Ball_Y_Step;
						  
					  else if ( (Ball_X_Pos + Ball_Size) >= Ball_X_Max )  // Ball is at the Right edge, BOUNCE!
					  begin  Ball_X_Motion <= (~ (Ball_X_Step) + 1'b1);  // 2's complement.
//						  Ball_Y_Pos <= Ball_Y_Center;
//						  Ball_X_Pos <= Ball_X_Center;
//						  Ball_X_Motion <= 3;
//						  Ball_Y_Motion <= -3;
						  Score1 <= (Score1+1'b1);
					  end	  
					 else if ( (Ball_X_Pos - Ball_Size) <= Ball_X_Min)
					 begin// Ball is at the Left edge, BOUNCE!
//						  Ball_Y_Pos <= Ball_Y_Center;
//						  Ball_X_Pos <= Ball_X_Center;
//						  Ball_X_Motion <= -3;
//						  Ball_Y_Motion <= 3;
						  Ball_X_Motion <= (Ball_X_Step);
						  Score2 <= (Score2+1'b1);
					 end	  
					 else 
						  Ball_Y_Motion <= Ball_Y_Motion;  // Ball is somewhere in the middle, don't bounce, just keep moving
						  
					 
					 Ball_Y_Pos <= (Ball_Y_Pos + Ball_Y_Motion);  // Update ball position
					 Ball_X_Pos <= (Ball_X_Pos + Ball_X_Motion);
				 end 
				 else begin
					 Ball_Y_Pos <= Ball_Y_Center;
					 Ball_X_Pos <= Ball_X_Center;
				 end	 
		end  
    end
       
    assign BallX = Ball_X_Pos;
   
    assign BallY = Ball_Y_Pos;
   
    assign BallS = Ball_Size;
    

endmodule